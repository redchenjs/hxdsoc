/*
 * exu2mem.sv
 *
 *  Created on: 2021-05-29 22:01
 *      Author: Jack Chen <redchenjs@live.com>
 */

module exu2mem #(
    parameter XLEN = 32
) (
    input logic clk_i,
    input logic rst_n_i
);

endmodule
