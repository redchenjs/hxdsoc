/*
 * config.sv
 *
 *  Created on: 2021-08-18 19:51
 *      Author: Jack Chen <redchenjs@live.com>
 */

`ifndef _CONFIG_SV_
`define _CONFIG_SV_

/* Base ISA */
`define CONFIG_ISA_RV32I

/* Extensions */
`define CONFIG_ISA_RV32C

`endif
