/*
 * config.sv
 *
 *  Created on: 2021-05-20 16:11
 *      Author: Jack Chen <redchenjs@live.com>
 */

parameter XLEN = 32;
