/*
 * mem2wb.sv
 *
 *  Created on: 2021-05-29 22:01
 *      Author: Jack Chen <redchenjs@live.com>
 */

module mem2wb #(
    parameter XLEN = 32
) (
    input logic clk_i,
    input logic rst_n_i
);

endmodule
